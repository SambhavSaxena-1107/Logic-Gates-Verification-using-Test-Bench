module nand_design(
    input wire A,
    input wire B,
    output wire Y
);
    assign Y = ~(A & B);
endmodule



