module not_design(
    input wire A,
    output wire Y
);
    assign Y = ~A ;
endmodule

